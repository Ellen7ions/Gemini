`timescale 1ns / 1ps

module ifu_2 (
    
);
    
endmodule