`timescale 1ns / 1ps

module ifu_1 (
    
);

endmodule