`timescale 1ns / 1ps

module ex (
    input   wire    clk,
    input   wire    rst,
    
    // control signals

    // data signals

    // output
);

endmodule