`timescale 1ns / 1ps

module d_cache (
    
);

endmodule